`timescale 1ns/1ps 
module mackey_TB;

	reg clk, rst, start;
	reg [7:0] ix1, ix2, ix3, ix4, ix5, ix6, ix7, ix8, ix9, ix10;
	reg [7:0] ix11, ix12, ix13, ix14, ix15, ix16, ix17, ix18, ix19, ix20;
	reg [9:0] instrucao;
	reg flagInst;

	wire oFlagRede;
	wire [7:0] oR1, oR2, oR3, oR4, oR5, oR6, oR7, oR8, oR9, oR10;
	wire [7:0] oR11, oR12, oR13, oR14, oR15, oR16, oR17, oR18, oR19, oR20;

	
	redeGeral r(clk, rst, start,
					instrucao, 
					flagInst, 
					ix1, ix2, ix3, ix4, ix5, ix6, ix7, ix8, ix9, ix10, ix11, ix12, ix13, ix14, ix15, ix16, ix17, ix18, ix19, ix20, 
					oR1, oR2, oR3, oR4, oR5, oR6, oR7, oR8, oR9, oR10, oR11, oR12, oR13, oR14, oR15, oR16, oR17, oR18, oR19, oR20, 
					oFlagRede
					); 
				
initial 
begin
	clk = 1'b0;
	rst = 1'b0;
	start = 1'b1;
	flagInst = 1'b1;
	instrucao = 10'b00_00001_0_00;
		
	ix1 = 8'b00000000; ix2 = 8'b00011101;
			
	#20 rst = 1'b1; 
		
	#20 flagInst = 1'b0; // CAPTURA A PRIMEIRA INSTRUÇÃO
		
	#20 flagInst = 1'b1;
	instrucao = 10'b10_00011_1_11;
		
	#20 flagInst = 1'b0; // CAPTURA A SEGUNDA INSTRUÇÃO
		
	#20 flagInst = 1'b1;
	instrucao = 10'b11_00000_1_01;
		
	#20 flagInst = 1'b0; // CAPTURA A TERCEIRA INSTRUÇÃO
	#20 flagInst = 1'b1;

	#1300 start = 1'b0; ix1 = 8'b00011101; ix2 = 8'b00011101; #20 start = 1'b1;
	#1300 start = 1'b0; ix1 = 8'b00011101; ix2 = 8'b00011100; #20 start = 1'b1;
	#1300 start = 1'b0; ix1 = 8'b00011100; ix2 = 8'b00011100; #20 start = 1'b1;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00001111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001111; ix2 = 8'b00001111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001111; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00101001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101001; ix2 = 8'b00101001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101001; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00001111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001111; ix2 = 8'b00001110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001110; ix2 = 8'b00001101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001101; ix2 = 8'b00001101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001101; ix2 = 8'b00001101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001101; ix2 = 8'b00001110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001110; ix2 = 8'b00001111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001111; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00101001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101001; ix2 = 8'b00101001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101001; ix2 = 8'b00101001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101001; ix2 = 8'b00101001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101001; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00001111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001111; ix2 = 8'b00001110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001110; ix2 = 8'b00001101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001101; ix2 = 8'b00001100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001100; ix2 = 8'b00001100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001100; ix2 = 8'b00001101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001101; ix2 = 8'b00001110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001110; ix2 = 8'b00001111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001111; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00001111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001111; ix2 = 8'b00001110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001110; ix2 = 8'b00001110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001110; ix2 = 8'b00001110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001110; ix2 = 8'b00001111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001111; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00100000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100000; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011010; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00101001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101001; ix2 = 8'b00101001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101001; ix2 = 8'b00101010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101010; ix2 = 8'b00101010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101010; ix2 = 8'b00101010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101010; ix2 = 8'b00101010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101010; ix2 = 8'b00101010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101010; ix2 = 8'b00101001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101001; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010110; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010001; ix2 = 8'b00010000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010000; ix2 = 8'b00001111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001111; ix2 = 8'b00001110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001110; ix2 = 8'b00001101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001101; ix2 = 8'b00001100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001100; ix2 = 8'b00001100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001100; ix2 = 8'b00001100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001100; ix2 = 8'b00001100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001100; ix2 = 8'b00001101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001101; ix2 = 8'b00001111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00001111; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011110; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100011; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100101; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00101000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00101000; ix2 = 8'b00100111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100111; ix2 = 8'b00100110; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100110; ix2 = 8'b00100100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100100; ix2 = 8'b00100010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100010; ix2 = 8'b00100001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00100001; ix2 = 8'b00011111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011111; ix2 = 8'b00011101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011101; ix2 = 8'b00011100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011100; ix2 = 8'b00011011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011011; ix2 = 8'b00011001; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011001; ix2 = 8'b00011000; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00011000; ix2 = 8'b00010111; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010111; ix2 = 8'b00010101; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010101; ix2 = 8'b00010100; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010100; ix2 = 8'b00010011; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010011; ix2 = 8'b00010010; #20 start = 1'b0;
	#1300 start = 1'b1; ix1 = 8'b00010010; ix2 = 8'b00010001; #20 start = 1'b0;
	
	#1300 $stop;
end
	
	always
	begin
		#10 clk = 1'b1;
		#10 clk = 1'b0;
	end

	
endmodule

`timescale 1ns/1ps //valor de fundo/precisao
module iris_TB;

	reg clk, rst, start;
	
	reg [7:0] ix1, ix2, ix3, ix4, ix5, ix6, ix7, ix8, ix9, ix10;
	reg [7:0] ix11, ix12, ix13, ix14, ix15, ix16, ix17, ix18, ix19, ix20;
	
	reg [9:0] instrucao;
	reg flagInst;
	
	wire oFlagRede;
	wire [7:0] oR1, oR2, oR3, oR4, oR5, oR6, oR7, oR8, oR9, oR10;
	wire [7:0] oR11, oR12, oR13, oR14, oR15, oR16, oR17, oR18, oR19, oR20;
	
	redeGeral r(clk, rst, start, 
					instrucao, 
					flagInst, 
					ix1, ix2, ix3, ix4, ix5, ix6, ix7, ix8, ix9, ix10, ix11, ix12, ix13, ix14, ix15, ix16, ix17, ix18, ix19, ix20,
					oR1, oR2, oR3, oR4, oR5, oR6, oR7, oR8, oR9, oR10, oR11, oR12, oR13, oR14, oR15, oR16, oR17, oR18, oR19, oR20,
					oFlagRede
					); 
				
initial 
begin	
		clk = 1'b0;
		rst = 1'b0;
		start = 1'b1;
		flagInst = 1'b1;
		instrucao = 10'b00_00011_0_00;
		
		ix1 = 8'b00011100; ix2 = 8'b01001111; ix3 = 8'b00001000; ix4 = 8'b00000101;
				
		#50 rst = 1'b1; 
		
		#120 flagInst = 1'b0; // CAPTURA A PRIMEIRA INSTRUÇÃO
		
		#40 flagInst = 1'b1;
		instrucao = 10'b10_00111_1_11;
		
		#40 flagInst = 1'b0; // CAPTURA A SEGUNDA INSTRUÇÃO
		
		#40 flagInst = 1'b1;
		instrucao = 10'b10_00010_1_11;
		
		#40 flagInst = 1'b0; // CAPTURA A TERCEIRA INSTRUÇÃO
		
		#40 flagInst = 1'b1;
		#40 instrucao = 10'b11_00010_1_01;
		
		#40 flagInst = 1'b0; // CAPTURA A QUARTA INSTRUÇÃO
		#40 flagInst = 1'b1;
		
		
		#10000 start = 1'b0; ix1 = 8'b00010101; ix2 = 8'b00110100; ix3 = 8'b00001000; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00001110; ix2 = 8'b00111111; ix3 = 8'b00000110; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00001010; ix2 = 8'b00111010; ix3 = 8'b00001010; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011000; ix2 = 8'b01010100; ix3 = 8'b00001000; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00100110; ix2 = 8'b01100100; ix3 = 8'b00001111; ix4 = 8'b00001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00001010; ix2 = 8'b01001010; ix3 = 8'b00001000; ix4 = 8'b00001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011000; ix2 = 8'b01001010; ix3 = 8'b00001010; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00000011; ix2 = 8'b00101111; ix3 = 8'b00001000; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00010101; ix2 = 8'b00111010; ix3 = 8'b00001010; ix4 = 8'b00000000; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00100110; ix2 = 8'b01011001; ix3 = 8'b00001010; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00010001; ix2 = 8'b01001010; ix3 = 8'b00001100; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00010001; ix2 = 8'b00110100; ix3 = 8'b00001000; ix4 = 8'b00000000; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00000000; ix2 = 8'b00110100; ix3 = 8'b00000010; ix4 = 8'b00000000; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110100; ix2 = 8'b01101001; ix3 = 8'b00000100; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110001; ix2 = 8'b01111111; ix3 = 8'b00001010; ix4 = 8'b00001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00100110; ix2 = 8'b01100100; ix3 = 8'b00000110; ix4 = 8'b00001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011100; ix2 = 8'b01001111; ix3 = 8'b00001000; ix4 = 8'b00001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110001; ix2 = 8'b01011111; ix3 = 8'b00001111; ix4 = 8'b00001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011100; ix2 = 8'b01011111; ix3 = 8'b00001010; ix4 = 8'b00001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00100110; ix2 = 8'b01001010; ix3 = 8'b00001111; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011100; ix2 = 8'b01011001; ix3 = 8'b00001010; ix4 = 8'b00001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00001010; ix2 = 8'b01010100; ix3 = 8'b00000000; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011100; ix2 = 8'b01000100; ix3 = 8'b00001111; ix4 = 8'b00010101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00010001; ix2 = 8'b01001010; ix3 = 8'b00010011; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011000; ix2 = 8'b00110100; ix3 = 8'b00001100; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011000; ix2 = 8'b01001010; ix3 = 8'b00001100; ix4 = 8'b00001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011111; ix2 = 8'b01001111; ix3 = 8'b00001010; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011111; ix2 = 8'b01001010; ix3 = 8'b00001000; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00001110; ix2 = 8'b00111111; ix3 = 8'b00001100; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00010001; ix2 = 8'b00111010; ix3 = 8'b00001100; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00100110; ix2 = 8'b01001010; ix3 = 8'b00001010; ix4 = 8'b00001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011111; ix2 = 8'b01101111; ix3 = 8'b00001010; ix4 = 8'b00000000; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101010; ix2 = 8'b01110100; ix3 = 8'b00001000; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00010101; ix2 = 8'b00111010; ix3 = 8'b00001010; ix4 = 8'b00000000; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011000; ix2 = 8'b00111111; ix3 = 8'b00000100; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101010; ix2 = 8'b01001111; ix3 = 8'b00000110; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00010101; ix2 = 8'b00111010; ix3 = 8'b00001010; ix4 = 8'b00000000; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00000011; ix2 = 8'b00110100; ix3 = 8'b00000110; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011100; ix2 = 8'b01001010; ix3 = 8'b00001010; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011000; ix2 = 8'b01001111; ix3 = 8'b00000110; ix4 = 8'b00001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00000111; ix2 = 8'b00001111; ix3 = 8'b00000110; ix4 = 8'b00001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00000011; ix2 = 8'b00111111; ix3 = 8'b00000110; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011000; ix2 = 8'b01001111; ix3 = 8'b00001100; ix4 = 8'b00011010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011100; ix2 = 8'b01011111; ix3 = 8'b00010011; ix4 = 8'b00001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00010001; ix2 = 8'b00110100; ix3 = 8'b00001000; ix4 = 8'b00001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011100; ix2 = 8'b01011111; ix3 = 8'b00001100; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00001010; ix2 = 8'b00111111; ix3 = 8'b00001000; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00100011; ix2 = 8'b01011001; ix3 = 8'b00001010; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011000; ix2 = 8'b01000100; ix3 = 8'b00001000; ix4 = 8'b00000101; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01011111; ix2 = 8'b00111111; ix3 = 8'b01001111; ix4 = 8'b01000100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001010; ix2 = 8'b00111111; ix3 = 8'b01001011; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01011011; ix2 = 8'b00111010; ix3 = 8'b01010011; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101010; ix2 = 8'b00001111; ix3 = 8'b01000000; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001101; ix2 = 8'b00101010; ix3 = 8'b01001101; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110001; ix2 = 8'b00101010; ix3 = 8'b01001011; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000110; ix2 = 8'b01000100; ix3 = 8'b01001111; ix4 = 8'b01001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00010101; ix2 = 8'b00010101; ix3 = 8'b00110001; ix4 = 8'b00101111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01010001; ix2 = 8'b00101111; ix3 = 8'b01001101; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011111; ix2 = 8'b00100101; ix3 = 8'b00111110; ix4 = 8'b01000100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011000; ix2 = 8'b00000000; ix3 = 8'b00110101; ix4 = 8'b00101111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111000; ix2 = 8'b00110100; ix3 = 8'b01000100; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111011; ix2 = 8'b00001010; ix3 = 8'b01000000; ix4 = 8'b00101111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111111; ix2 = 8'b00101111; ix3 = 8'b01001111; ix4 = 8'b01000100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101101; ix2 = 8'b00101111; ix3 = 8'b00110111; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01010100; ix2 = 8'b00111010; ix3 = 8'b01001001; ix4 = 8'b01000100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101101; ix2 = 8'b00110100; ix3 = 8'b01001011; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110100; ix2 = 8'b00100101; ix3 = 8'b01000010; ix4 = 8'b00101111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000011; ix2 = 8'b00001010; ix3 = 8'b01001011; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101101; ix2 = 8'b00011010; ix3 = 8'b00111110; ix4 = 8'b00110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111000; ix2 = 8'b00111111; ix3 = 8'b01010001; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111111; ix2 = 8'b00101010; ix3 = 8'b01000000; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000110; ix2 = 8'b00011010; ix3 = 8'b01010011; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111111; ix2 = 8'b00101010; ix3 = 8'b01001111; ix4 = 8'b00111010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001010; ix2 = 8'b00101111; ix3 = 8'b01000111; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01010001; ix2 = 8'b00110100; ix3 = 8'b01001001; ix4 = 8'b01000100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01011000; ix2 = 8'b00101010; ix3 = 8'b01010001; ix4 = 8'b01000100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01010100; ix2 = 8'b00110100; ix3 = 8'b01010110; ix4 = 8'b01010100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111011; ix2 = 8'b00101111; ix3 = 8'b01001011; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110001; ix2 = 8'b00011111; ix3 = 8'b00110101; ix4 = 8'b00101111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101010; ix2 = 8'b00010101; ix3 = 8'b00111100; ix4 = 8'b00110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101010; ix2 = 8'b00010101; ix3 = 8'b00111010; ix4 = 8'b00101111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110100; ix2 = 8'b00100101; ix3 = 8'b00111110; ix4 = 8'b00111010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111011; ix2 = 8'b00100101; ix3 = 8'b01011000; ix4 = 8'b01001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00100110; ix2 = 8'b00110100; ix3 = 8'b01001011; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111011; ix2 = 8'b01001010; ix3 = 8'b01001011; ix4 = 8'b01001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01010100; ix2 = 8'b00111010; ix3 = 8'b01001111; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000110; ix2 = 8'b00001111; ix3 = 8'b01001001; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101101; ix2 = 8'b00110100; ix3 = 8'b01000010; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101010; ix2 = 8'b00011010; ix3 = 8'b01000000; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101010; ix2 = 8'b00011111; ix3 = 8'b01001001; ix4 = 8'b00111010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111111; ix2 = 8'b00110100; ix3 = 8'b01001101; ix4 = 8'b01000100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110100; ix2 = 8'b00011111; ix3 = 8'b01000000; ix4 = 8'b00111010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011000; ix2 = 8'b00001111; ix3 = 8'b00110001; ix4 = 8'b00101111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101101; ix2 = 8'b00100101; ix3 = 8'b01000100; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110001; ix2 = 8'b00110100; ix3 = 8'b01000100; ix4 = 8'b00111010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110001; ix2 = 8'b00101111; ix3 = 8'b01000100; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000011; ix2 = 8'b00101111; ix3 = 8'b01000111; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00011100; ix2 = 8'b00011010; ix3 = 8'b00101011; ix4 = 8'b00110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110001; ix2 = 8'b00101010; ix3 = 8'b01000010; ix4 = 8'b00111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000110; ix2 = 8'b01000100; ix3 = 8'b01101011; ix4 = 8'b01111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110100; ix2 = 8'b00100101; ix3 = 8'b01011000; ix4 = 8'b01011111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01100010; ix2 = 8'b00110100; ix3 = 8'b01101001; ix4 = 8'b01101001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000110; ix2 = 8'b00101111; ix3 = 8'b01100011; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001101; ix2 = 8'b00110100; ix3 = 8'b01100111; ix4 = 8'b01101111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01110100; ix2 = 8'b00110100; ix3 = 8'b01111000; ix4 = 8'b01101001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00010101; ix2 = 8'b00011010; ix3 = 8'b01001011; ix4 = 8'b01010100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01101001; ix2 = 8'b00101111; ix3 = 8'b01110010; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01010100; ix2 = 8'b00011010; ix3 = 8'b01100111; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01100110; ix2 = 8'b01010100; ix3 = 8'b01101101; ix4 = 8'b01111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001101; ix2 = 8'b00111111; ix3 = 8'b01011000; ix4 = 8'b01100100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001010; ix2 = 8'b00100101; ix3 = 8'b01011100; ix4 = 8'b01011111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01011000; ix2 = 8'b00110100; ix3 = 8'b01100000; ix4 = 8'b01101001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110001; ix2 = 8'b00011010; ix3 = 8'b01010110; ix4 = 8'b01100100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110100; ix2 = 8'b00101010; ix3 = 8'b01011000; ix4 = 8'b01111001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001010; ix2 = 8'b00111111; ix3 = 8'b01011100; ix4 = 8'b01110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001101; ix2 = 8'b00110100; ix3 = 8'b01100000; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01110111; ix2 = 8'b01011111; ix3 = 8'b01111010; ix4 = 8'b01101111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01110111; ix2 = 8'b00011111; ix3 = 8'b01111111; ix4 = 8'b01110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111011; ix2 = 8'b00001010; ix3 = 8'b01010110; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01011011; ix2 = 8'b00111111; ix3 = 8'b01100101; ix4 = 8'b01110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00101101; ix2 = 8'b00101010; ix3 = 8'b01010011; ix4 = 8'b01100100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01110111; ix2 = 8'b00101010; ix3 = 8'b01111010; ix4 = 8'b01100100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000110; ix2 = 8'b00100101; ix3 = 8'b01010011; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01010100; ix2 = 8'b01000100; ix3 = 8'b01100101; ix4 = 8'b01101001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01100110; ix2 = 8'b00111111; ix3 = 8'b01101011; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000011; ix2 = 8'b00101010; ix3 = 8'b01010001; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111111; ix2 = 8'b00110100; ix3 = 8'b01010011; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001010; ix2 = 8'b00101010; ix3 = 8'b01100011; ix4 = 8'b01101001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01100110; ix2 = 8'b00110100; ix3 = 8'b01100111; ix4 = 8'b01001111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01101101; ix2 = 8'b00101010; ix3 = 8'b01101101; ix4 = 8'b01011111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01111111; ix2 = 8'b01011111; ix3 = 8'b01110100; ix4 = 8'b01100100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001010; ix2 = 8'b00101010; ix3 = 8'b01100011; ix4 = 8'b01101111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000110; ix2 = 8'b00101010; ix3 = 8'b01011000; ix4 = 8'b01001010; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111111; ix2 = 8'b00011111; ix3 = 8'b01100011; ix4 = 8'b01000100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01110111; ix2 = 8'b00110100; ix3 = 8'b01101101; ix4 = 8'b01110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000110; ix2 = 8'b01001010; ix3 = 8'b01100011; ix4 = 8'b01111001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001010; ix2 = 8'b00111010; ix3 = 8'b01100000; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111011; ix2 = 8'b00110100; ix3 = 8'b01010001; ix4 = 8'b01011001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01011011; ix2 = 8'b00111010; ix3 = 8'b01011110; ix4 = 8'b01101001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01010100; ix2 = 8'b00111010; ix3 = 8'b01100011; ix4 = 8'b01111001; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01011011; ix2 = 8'b00111010; ix3 = 8'b01011000; ix4 = 8'b01110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00110100; ix2 = 8'b00100101; ix3 = 8'b01011000; ix4 = 8'b01011111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01011000; ix2 = 8'b00111111; ix3 = 8'b01101001; ix4 = 8'b01110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01010100; ix2 = 8'b01000100; ix3 = 8'b01100101; ix4 = 8'b01111111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01010100; ix2 = 8'b00110100; ix3 = 8'b01011010; ix4 = 8'b01110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000110; ix2 = 8'b00011010; ix3 = 8'b01010110; ix4 = 8'b01011111; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01001101; ix2 = 8'b00110100; ix3 = 8'b01011010; ix4 = 8'b01100100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b01000011; ix2 = 8'b01001010; ix3 = 8'b01011110; ix4 = 8'b01110100; #40 start = 1'b1;
		#10000 start = 1'b0; ix1 = 8'b00111000; ix2 = 8'b00110100; ix3 = 8'b01011000; ix4 = 8'b01011001; #40 start = 1'b1;


		#20000 $stop;
end
	
	always
	begin
		#20 clk = 1'b1;
		#20 clk = 1'b0;
	end

	
endmodule

module unidadeMemoria(clk, rst,     // CLOCK E RESET DO SISTEMA
							 iStartCarga,  // FLAG DE INICIO DA BUSCA DOS DADOS NAS MEMORIAS
							 iFlagCamada,   // INDICA QUE A CAMADA INICIOU SUA EXECUÇÃO
							 iCamada,      // NUMERO DA CAMADA QUE ESTA' EM EXECUCAO
							 iQtdEntradas,       // QUANTIDADE DE ENTRADAS DA CAMADA
							 iQtdNeuro,    // QUANTIDADE DE NEURONIOS DA CAMADA
							 oW,           // PESOS DAS ENTRADAS
							 oBias,        // BIAS DOS NEURONIOS
							 oPesosOK);    // FLAG DE SAIDA DO CARREGAMENTO
	
	input clk, rst;
	input iStartCarga, iFlagCamada;
	input [1:0] iCamada;
	input [4:0] iQtdEntradas, iQtdNeuro;
	
	output reg [15:0] oW [0:399]; 
	output reg oPesosOK; 
	output reg [15:0] oBias [0:19];

	reg [5:0] i; // CONTAGEM DE NEURONIOS
	reg [6:0] addr; // ENDERECO 
	reg flagLeitura, flagMemoria; // HABILITAM AS MEMORIAS
	wire [15:0] oS1, oS2, oS3, oS4, oS5, oS6, oS7, oS8, oS9, oS10, oS11, oS12, oS13, oS14, oS15, oS16, oS17, oS18, oS19, oS20, oSBias; // SAIDAS AUXILIARES DAS MEMORIAS
	
	(* syn_encoding = "safe" *) reg [1:0] atual;  
	parameter S0 = 2'b00, S1 = 2'b01, S2 = 2'b10, S3 = 2'b11; // ESTADOS

	memoria_neuro1 m1(clk, addr, oS1, flagLeitura, flagMemoria);
	memoria_neuro2 m2(clk, addr, oS2, flagLeitura, flagMemoria);
	memoria_neuro3 m3(clk, addr, oS3, flagLeitura, flagMemoria);
	memoria_neuro4 m4(clk, addr, oS4, flagLeitura, flagMemoria);
	memoria_neuro5 m5(clk, addr, oS5, flagLeitura, flagMemoria);
	memoria_neuro6 m6(clk, addr, oS6, flagLeitura, flagMemoria);
	memoria_neuro7 m7(clk, addr, oS7, flagLeitura, flagMemoria);
	memoria_neuro8 m8(clk, addr, oS8, flagLeitura, flagMemoria);
	memoria_neuro9 m9(clk, addr, oS9, flagLeitura, flagMemoria);
	memoria_neuro10 m10(clk, addr, oS10, flagLeitura, flagMemoria);
	memoria_neuro11 m11(clk, addr, oS11, flagLeitura, flagMemoria);
	memoria_neuro12 m12(clk, addr, oS12, flagLeitura, flagMemoria);
	memoria_neuro13 m13(clk, addr, oS13, flagLeitura, flagMemoria);
	memoria_neuro14 m14(clk, addr, oS14, flagLeitura, flagMemoria);
	memoria_neuro15 m15(clk, addr, oS15, flagLeitura, flagMemoria);
	memoria_neuro16 m16(clk, addr, oS16, flagLeitura, flagMemoria);
	memoria_neuro17 m17(clk, addr, oS17, flagLeitura, flagMemoria);
	memoria_neuro18 m18(clk, addr, oS18, flagLeitura, flagMemoria);
	memoria_neuro19 m19(clk, addr, oS19, flagLeitura, flagMemoria);
	memoria_neuro20 m20(clk, addr, oS20, flagLeitura, flagMemoria);
	
	memoria_bias m21(clk, addr, oSBias, flagLeitura, flagMemoria);

   always @(negedge clk, negedge rst)
	begin
		if(~rst)
		begin
			oPesosOK = 1'b0;
			// ZERAR PESOS E BIAS
			oW = '{{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
					 {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}};
					 
			oBias = '{{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}},
						{16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}, {16{1'b0}}};
						
			atual <= S0;
		end
		else
			case (atual) 
				S0: // PREPARA A BUSCA - ZERA OS FLAGS DE CONTROLE
				begin
					oPesosOK = 1'b0;
					i = 6'b000000;
					flagLeitura = 1'b0;
					flagMemoria = 1'b0;
					if(iStartCarga)
						atual <= S1;
					else
						atual <= S0;
				end
				S1: // INICIA A BUSCA - CALCULA O ENDERECO
				begin
			      oPesosOK = 1'b0;
					addr = {iCamada,i[4:0]};	
					flagLeitura = 1'b1;
					flagMemoria = 1'b1;
					atual <= S2;
				end
				S2: // ENCERRA A BUSCA - RECEBE OS RESULTADOS
				begin
					oPesosOK = 1'b0;
					oW[9'b000000000 + i[4:0]] = oS1;
					oW[9'b000010100 + i[4:0]] = oS2;
					oW[9'b000101000 + i[4:0]] = oS3;
					oW[9'b000111100 + i[4:0]] = oS4;
					oW[9'b001010000 + i[4:0]] = oS5;
					oW[9'b001100100 + i[4:0]] = oS6;
					oW[9'b001111000 + i[4:0]] = oS7;
					oW[9'b010001100 + i[4:0]] = oS8;
					oW[9'b010100000 + i[4:0]] = oS9;
					oW[9'b010110100 + i[4:0]] = oS10;
					oW[9'b011001000 + i[4:0]] = oS11;
					oW[9'b011011100 + i[4:0]] = oS12;
					oW[9'b011110000 + i[4:0]] = oS13;
					oW[9'b100000100 + i[4:0]] = oS14;
					oW[9'b100011000 + i[4:0]] = oS15;
					oW[9'b100101100 + i[4:0]] = oS16;
					oW[9'b101000000 + i[4:0]] = oS17;
					oW[9'b101010100 + i[4:0]] = oS18;
					oW[9'b101101000 + i[4:0]] = oS19;
					oW[9'b101111100 + i[4:0]] = oS20;
					
					oBias[i[4:0]] = oSBias;
					flagLeitura = 1'b0;
					flagMemoria = 1'b0;
					i = i + 6'b000001;
					if(i <= iQtdEntradas | i <= iQtdNeuro) // VERIFICA SE ACABOU
						atual <= S1;
					else
						atual <= S3;
				end
				S3: // ENCERRA O BLOCO
				begin
					oPesosOK = 1'b1;
					flagLeitura = 1'b0;
					flagMemoria = 1'b0;
					i = 6'b000000;
					if(iStartCarga | iFlagCamada)
					begin
						oPesosOK = 1'b0;
						atual <= S1;
					end
					else
						atual <= S3;
				end
			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 1
module memoria_neuro1(clk, iAddr, oS, iFlagLeitura, iFlagMem);
	input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0000111110011100; // CAMADA 1
				7'b0000001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0000000001000010; // CAMADA 2
				7'b0100001: oS <= 16'b1111111111011110; // CAMADA 2
				7'b0100010: oS <= 16'b0000000010010010; // CAMADA 2
				7'b0100011: oS <= 16'b0000000101100010; // CAMADA 2
				7'b0100100: oS <= 16'b1111111111111001; // CAMADA 2
				7'b0100101: oS <= 16'b0000000110100111; // CAMADA 2
				7'b0100110: oS <= 16'b0000001010010001; // CAMADA 2
				7'b0100111: oS <= 16'b0000010010111001; // CAMADA 2
				7'b0101000: oS <= 16'b1111111110110001; // CAMADA 2
				7'b0101001: oS <= 16'b1111111010010111; // CAMADA 2
				7'b0101010: oS <= 16'b1111111110011111; // CAMADA 2
				7'b0101011: oS <= 16'b0000000000110000; // CAMADA 2
				7'b0101100: oS <= 16'b1111111110111010; // CAMADA 2
				7'b0101101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 2
module memoria_neuro2(clk, iAddr, oS, iFlagLeitura, iFlagMem);
	input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0001000100011001; // CAMADA 1
				7'b0000001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0010100000000000; // CAMADA 2
				7'b0100001: oS <= 16'b1101100000000000; // CAMADA 2
				7'b0100010: oS <= 16'b0000011000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0100100: oS <= 16'b0000101000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0100111: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0101000: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0101010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101011: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0110010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4
			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 3
module memoria_neuro3(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b1111011000001110; // CAMADA 1
				7'b0000001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0001010000000000; // CAMADA 2
				7'b0100001: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0100010: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0000101000000000; // CAMADA 2
				7'b0100100: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0100101: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0100111: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101000: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101010: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110000: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000001000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4
			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 4
module memoria_neuro4(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0000011100110101; // CAMADA 1
				7'b0000001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0010100000000000; // CAMADA 2
				7'b0100001: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0100010: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0100011: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0100101: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100111: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101001: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101101: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101110: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000001000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0110001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000011000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 5
module memoria_neuro5(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0001010011000001; // CAMADA 1
				7'b0000001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0100001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100010: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100100: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0100110: oS <= 16'b0000101000000000; // CAMADA 2
				7'b0100111: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101000: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000001000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000011000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000101000000000; // CAMADA 2
				7'b0101111: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0110000: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0110010: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0111001: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0111010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000001000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000011000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000100000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 6
module memoria_neuro6(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b1111100000101111; // CAMADA 1
				7'b0000001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0100001: oS <= 16'b0001011000000000; // CAMADA 2
				7'b0100010: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0100101: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0100111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101001: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101010: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101100: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101101: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000001000000000; // CAMADA 2
				7'b0101111: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000101000000000; // CAMADA 2
				7'b0110011: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 7
module memoria_neuro7(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b1111100101000101; // CAMADA 1
				7'b0000001: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000010: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000100: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0000101: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000110: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0001001: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000110000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000011000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000101000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000110000000000; // CAMADA 1
				7'b0010000: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0010001: oS <= 16'b1111011000000000; // CAMADA 1
				7'b0010010: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0100001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100010: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0100101: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0100111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000011000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000101000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0110000: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0110010: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 8
module memoria_neuro8(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0000010101001011; // CAMADA 1
				7'b0000001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0000011: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000110000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000011000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000101000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000110000000000; // CAMADA 1
				7'b0001010: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0001011: oS <= 16'b1111011000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0001110: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001111: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010001: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0010010: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b1110110000000000; // CAMADA 2
				7'b0100001: oS <= 16'b0001010000000000; // CAMADA 2
				7'b0100010: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0100011: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0100100: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0100110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100111: oS <= 16'b0000011000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000101000000000; // CAMADA 2
				7'b0101001: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0101010: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0101011: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101101: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0101110: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101111: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0110010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 9
module memoria_neuro9(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0000101110110110; // CAMADA 1
				7'b0000001: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0000010: oS <= 16'b1111011000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000100: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0000101: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000110: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0001001: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001100: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0001101: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000001000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000101000000000; // CAMADA 1
				7'b0010001: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0010010: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0010011: oS <= 16'b1111011000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0001100000000000; // CAMADA 2
				7'b0100001: oS <= 16'b1110100000000000; // CAMADA 2
				7'b0100010: oS <= 16'b0001010000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0001000000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0100101: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0100111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101000: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101100: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101101: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000001000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000101000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0110010: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0110011: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 10
module memoria_neuro10(clk, iAddr, oS, iFlagLeitura, iFlagMem);
	input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0000011110001001; // CAMADA 1
				7'b0000001: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0000100: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0000111: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0001000: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0001101: oS <= 16'b1111011000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0010000: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010001: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0001010000000000; // CAMADA 2
				7'b0100001: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0100010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100011: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100110: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0100111: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101000: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101001: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101100: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0101101: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101111: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0110000: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 11
module memoria_neuro11(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b1111001110000010; // CAMADA 1
				7'b0000001: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0000010: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0000111: oS <= 16'b1111011000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0001010: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0001111: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0010010: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0001010000000000; // CAMADA 2
				7'b0100001: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0100010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0100100: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0100111: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0101010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101100: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101110: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0101111: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110001: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110010: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 12
module memoria_neuro12(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0001000001001100; // CAMADA 1
				7'b0000001: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0000100: oS <= 16'b1111011000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0000111: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001011: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0001100: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0001010000000000; // CAMADA 2
				7'b0100001: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0100010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100011: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0100111: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101011: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0101100: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0110001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110010: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 13
module memoria_neuro13(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0000111011110000; // CAMADA 1
				7'b0000001: oS <= 16'b1111011000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0000100: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0001001: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0001101: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0010000: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b1110100000000000; // CAMADA 2
				7'b0100001: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0100010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100011: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0100111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101000: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101101: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101111: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0110000: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 14
module memoria_neuro14(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0000110000000000; // CAMADA 1
				7'b0000001: oS <= 16'b1111101000000000; // CAMADA 1
				7'b0000010: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000011: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0000111: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001001: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0001010: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001011: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001110: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0001111: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000001000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0010010: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000110000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0001100000000000; // CAMADA 2
				7'b0100001: oS <= 16'b1111101000000000; // CAMADA 2
				7'b0100010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100011: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0100100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0100110: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0100111: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101011: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101110: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101111: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000001000000000; // CAMADA 2
				7'b0110001: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 15
module memoria_neuro15(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0000001: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0000010: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0000100: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0000101: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000110: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001001: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0001010: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0010000: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000110000000000; // CAMADA 1
				7'b0010011: oS <= 16'b1111000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0100001: oS <= 16'b0001000000000000; // CAMADA 2
				7'b0100010: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0100101: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101100: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0110000: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0110001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0110011: oS <= 16'b1111000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 16
module memoria_neuro16(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0000011: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0000100: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001010: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001110: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0010000: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0010001: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010010: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010011: oS <= 16'b1111011000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b1110110000000000; // CAMADA 2
				7'b0100001: oS <= 16'b0001010000000000; // CAMADA 2
				7'b0100010: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0100011: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101010: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101110: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110000: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110011: oS <= 16'b1111011000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4
			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 17
module memoria_neuro17(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0000001: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000111: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001110: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0001111: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010000: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000110000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b1111000000000000; // CAMADA 2
				7'b0100001: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0100010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100011: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100111: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101001: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101100: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101110: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0101111: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110000: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 18
module memoria_neuro18(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000001: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000100: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000101: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000111: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001001: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001110: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0010000: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0010001: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0100001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100101: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0100110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100111: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101001: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101110: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110000: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 19
module memoria_neuro19(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0000001: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000011: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000111: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0001000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001011: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0010000: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0010001: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b1111000000000000; // CAMADA 2
				7'b0100001: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0100010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100011: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100110: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100111: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101001: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101011: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110000: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0110001: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule

// MEMÓRIA PESOS NEURÔNIO 20
module memoria_neuro20(clk, iAddr, oS, iFlagLeitura, iFlagMem);
	input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0000001: oS <= 16'b1111100000000000; // CAMADA 1
				7'b0000010: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000100: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0000101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0000111: oS <= 16'b1111110000000000; // CAMADA 1
				7'b0001000: oS <= 16'b1111111000000000; // CAMADA 1
				7'b0001001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001010: oS <= 16'b0000010000000000; // CAMADA 1
				7'b0001011: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001101: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0001110: oS <= 16'b1111010000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000100000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000110000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0000011000000000; // CAMADA 2
				7'b0100001: oS <= 16'b1111100000000000; // CAMADA 2
				7'b0100010: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100100: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100111: oS <= 16'b1111110000000000; // CAMADA 2
				7'b0101000: oS <= 16'b1111111000000000; // CAMADA 2
				7'b0101001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000010000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0101110: oS <= 16'b1111010000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000100000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000110000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4
			endcase
	end
endmodule

// MEMÓRIA DO BIAS
module memoria_bias(clk, iAddr, oS, iFlagLeitura, iFlagMem);
input [6:0] iAddr;
	input iFlagLeitura;
	input iFlagMem;
	input clk;
	output reg [15:0] oS;

	always @ (posedge clk)
	begin
		if (iFlagLeitura | iFlagMem)
			case (iAddr)
				7'b0000000: oS <= 16'b1100010001000111; // CAMADA 1
				7'b0000001: oS <= 16'b1100101010010010; // CAMADA 1
				7'b0000010: oS <= 16'b0001101110001111; // CAMADA 1
				7'b0000011: oS <= 16'b1111001010111001; // CAMADA 1
				7'b0000100: oS <= 16'b1110011110011010; // CAMADA 1
				7'b0000101: oS <= 16'b0000011010010011; // CAMADA 1
				7'b0000110: oS <= 16'b0000001010011100; // CAMADA 1
				7'b0000111: oS <= 16'b0000001101010001; // CAMADA 1
				7'b0001000: oS <= 16'b0001011111100111; // CAMADA 1
				7'b0001001: oS <= 16'b0000110001110010; // CAMADA 1
				7'b0001010: oS <= 16'b1101110101001010; // CAMADA 1
				7'b0001011: oS <= 16'b0011001011111011; // CAMADA 1
				7'b0001100: oS <= 16'b0011100101110111; // CAMADA 1
				7'b0001101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0001111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0010111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011000: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011001: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011010: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011011: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011100: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011101: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011110: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0011111: oS <= 16'b0000000000000000; // CAMADA 1
				7'b0100000: oS <= 16'b0000000000011010; // CAMADA 2
				7'b0100001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0100111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0101111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0110111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111000: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111001: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111010: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111011: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111100: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111101: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111110: oS <= 16'b0000000000000000; // CAMADA 2
				7'b0111111: oS <= 16'b0000000000000000; // CAMADA 2
				7'b1000000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1000111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1001111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1010111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011000: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011001: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011010: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011011: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011100: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011101: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011110: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1011111: oS <= 16'b0000000000000000; // CAMADA 3
				7'b1100000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1100111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1101111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1110111: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111000: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111001: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111010: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111011: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111100: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111101: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111110: oS <= 16'b0000000000000000; // CAMADA 4
				7'b1111111: oS <= 16'b0000000000000000; // CAMADA 4

			endcase
	end
endmodule
